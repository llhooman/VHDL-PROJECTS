LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY carry_lookahead_adder IS
    PORT (
        A : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0):="1000011111001000";
        B : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0):="0000011111000001";
        CMINUS1 : INOUT STD_LOGIC:='0';
        S : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY carry_lookahead_adder;

ARCHITECTURE rtl OF carry_lookahead_adder IS
    SIGNAL C0, C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11, C12, C13, C14, C15 : STD_LOGIC;
    SIGNAL G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15 : STD_LOGIC;
    SIGNAL P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15 : STD_LOGIC;
BEGIN
    --Gi = Ai AND Bi
    G0 <= A(0) AND B(0);
    G1 <= A(1) AND B(1);
    G2 <= A(2) AND B(2);
    G3 <= A(3) AND B(3);
    G4 <= A(4) AND B(4);
    G5 <= A(5) AND B(5);
    G6 <= A(6) AND B(6);
    G7 <= A(7) AND B(7);
    G8 <= A(8) AND B(8);
    G9 <= A(9) AND B(9);
    G10 <= A(10) AND B(10);
    G11 <= A(11) AND B(11);
    G12 <= A(12) AND B(12);
    G13 <= A(13) AND B(13);
    G14 <= A(14) AND B(14);
    G15 <= A(15) AND B(15);
    --Pi = Ai XOR Bi
    P0 <= A(0) XOR B(0);
    P1 <= A(1) XOR B(1);
    P2 <= A(2) XOR B(2);
    P3 <= A(3) XOR B(3);
    P4 <= A(4) XOR B(4);
    P5 <= A(5) XOR B(5);
    P6 <= A(6) XOR B(6);
    P7 <= A(7) XOR B(7);
    P8 <= A(8) XOR B(8);
    P9 <= A(9) XOR B(9);
    P10 <= A(10) XOR B(10);
    P11 <= A(11) XOR B(11);
    P12 <= A(12) XOR B(12);
    P13 <= A(13) XOR B(13);
    P14 <= A(14) XOR B(14);
    P15 <= A(15) XOR B(15);

    --calculating the carries
    C0 <= G0 OR (P0 AND CMINUS1);
    C1 <= G1 OR (P1 AND G0) OR (P1 AND P0 AND CMINUS1);
    C2 <= G2 OR (P2 AND G1) OR (P2 AND P1 AND G0) OR (P2 AND P1 AND P0 AND CMINUS1);
    C3 <= G3 OR (P3 AND G2) OR (P3 AND P2 AND G1) OR (P3 AND P2 AND P1 AND G0) OR (P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C4 <= G4 OR (P4 AND G3) OR (P4 AND P3 AND G2) OR (P4 AND P3 AND P2 AND G1) OR (P4 AND P3 AND P2 AND P1 AND G0) OR (P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C5 <= G5 OR (P5 AND G4) OR (P5 AND P4 AND G3) OR (P5 AND P4 AND P3 AND G2) OR (P5 AND P4 AND P3 AND P2 AND G1) OR (P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C6 <= G6 OR (P6 AND G5) OR (P6 AND P5 AND G4) OR (P6 AND P5 AND P4 AND G3) OR (P6 AND P5 AND P4 AND P3 AND G2) OR (P6 AND P5 AND P4 AND P3 AND P2 AND G1) OR (P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C7 <= G7 OR (P7 AND G6) OR (P7 AND P6 AND G5) OR (P7 AND P6 AND P5 AND G4) OR (P7 AND P6 AND P5 AND P4 AND G3) OR (P7 AND P6 AND P5 AND P4 AND P3 AND G2) OR (P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND G1) OR (P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C8 <= G8 OR (P8 AND G7) OR (P8 AND P7 AND G6) OR (P8 AND P7 AND P6 AND G5) OR (P8 AND P7 AND P6 AND P5 AND G4) OR (P8 AND P7 AND P6 AND P5 AND P4 AND G3) OR (P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND G2) OR (P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND G1) OR (P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C9 <= G9 OR (P9 AND G8) OR (P9 AND P8 AND G7) OR (P9 AND P8 AND P7 AND G6) OR (P9 AND P8 AND P7 AND P6 AND G5) OR (P9 AND P8 AND P7 AND P6 AND P5 AND G4) OR (P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND G3) OR (P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND G2) OR (P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND G1) OR (P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C10 <= G10 OR (P10 AND G9) OR (P10 AND P9 AND G8) OR (P10 AND P9 AND P8 AND G7) OR (P10 AND P9 AND P8 AND P7 AND G6) OR (P10 AND P9 AND P8 AND P7 AND P6 AND G5) OR (P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND G4) OR (P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND G3) OR (P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND G2) OR (P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND G1) OR (P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C11 <= G11 OR (P11 AND G10) OR (P11 AND P10 AND G9) OR (P11 AND P10 AND P9 AND G8) OR (P11 AND P10 AND P9 AND P8 AND G7) OR (P11 AND P10 AND P9 AND P8 AND P7 AND G6) OR (P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND G5) OR (P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND G4) OR (P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND G3) OR (P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND G2) OR (P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND G1) OR (P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C12 <= G12 OR (P12 AND G11) OR (P12 AND P11 AND G10) OR (P12 AND P11 AND P10 AND G9) OR (P12 AND P11 AND P10 AND P9 AND G8) OR (P12 AND P11 AND P10 AND P9 AND P8 AND G7) OR (P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND G6) OR (P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND G5) OR (P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND G4) OR (P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND G3) OR (P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND G2) OR (P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND G1) OR (P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C13 <= G13 OR (P13 AND G12) OR (P13 AND P12 AND G11) OR (P13 AND P12 AND P11 AND G10) OR (P13 AND P12 AND P11 AND P10 AND G9) OR (P13 AND P12 AND P11 AND P10 AND P9 AND G8) OR (P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND G7) OR (P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND G6) OR (P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND G5) OR (P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND G4) OR (P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND G3) OR (P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND G2) OR (P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND G1) OR (P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C14 <= G14 OR (P14 AND G13) OR (P14 AND P13 AND G12) OR (P14 AND P13 AND P12 AND G11) OR (P14 AND P13 AND P12 AND P11 AND G10) OR (P14 AND P13 AND P12 AND P11 AND P10 AND G9) OR (P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND G8) OR (P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND G7) OR (P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND G6) OR (P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND G5) OR (P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND G4) OR (P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND G3) OR (P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND G2) OR (P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND G1) OR (P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);
    C15 <= G15 OR (P15 AND G14) OR (P15 AND P14 AND G13) OR (P15 AND P14 AND P13 AND G12) OR (P15 AND P14 AND P13 AND P12 AND G11) OR (P15 AND P14 AND P13 AND P12 AND P11 AND G10) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND G9) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND G8) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND G7) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND G6) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND G5) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND G4) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND G3) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND G2) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND G1) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND G0) OR (P15 AND P14 AND P13 AND P12 AND P11 AND P10 AND P9 AND P8 AND P7 AND P6 AND P5 AND P4 AND P3 AND P2 AND P1 AND P0 AND CMINUS1);

    --CALCULATING SUM
    S(0)<=A(0) XOR B(0) XOR CMINUS1;
    S(1)<=A(1) XOR B(1) XOR C0;
    S(2)<=A(2) XOR B(2) XOR C1;
    S(3)<=A(3) XOR B(3) XOR C2;
    S(4)<=A(4) XOR B(4) XOR C3;
    S(5)<=A(5) XOR B(5) XOR C4;
    S(6)<=A(6) XOR B(6) XOR C5;
    S(7)<=A(7) XOR B(7) XOR C6;
    S(8)<=A(8) XOR B(8) XOR C7;
    S(9)<=A(9) XOR B(9) XOR C8;
    S(10)<=A(10) XOR B(10) XOR C9;
    S(11)<=A(11) XOR B(11) XOR C10;
    S(12)<=A(12) XOR B(12) XOR C11;
    S(13)<=A(13) XOR B(13) XOR C12;
    S(14)<=A(14) XOR B(14) XOR C13;
    S(15)<=A(15) XOR B(15) XOR C14;
    
END ARCHITECTURE rtl;